`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2022/05/16 11:12:51
// Design Name: 
// Module Name: testbench
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module testbench();
reg                clk_in_p , clk_in_n;
reg       [3:0]    sw;                     //�ĸ����뿪�أ�������ʾ���ݵ�ת��
reg       [1:0]    key;                    //���������������ֱ��������ܵ�λѡ�����ֵĵ���
reg                rst;                    //ȫ�ָ�λ
wire      [7:0]    en;                     //�����ʹ���ź�
wire      [7:0]    disp1;                  //�����������ʾ
wire      [5:0]    led;
top top_sim(
    .clk_in_p(clk_in_p),
    .clk_in_n(clk_in_n),
    .rst(rst),
    .led(led),
    .sw(sw),
    .key(key),
    .en(en),
    .disp1(disp1)
);
initial    begin
    clk_in_p=0;
    clk_in_n=1;
    sw[3:0]=4'b0000;
    key[1:0]=2'b11;
    rst=1;
    #100000
    sw[3:0]=4'b0001;//�����յ�����
    #100000
    key[1:0]=2'b01;//���ǧλ��һ
    #10000000
    key[1:0]=2'b11;
    
    #100000
    sw[3:0]=4'b0011;//ʱ���������
    #100000
    key[1:0]=2'b01;//Сʱ��һ
    #10000000
    key[1:0]=2'b11;
//    #10000000
//    key[1:0]=2'b01;//Сʱ��һ
//    #10000000
//    key[1:0]=2'b11;
//    sw[3:0]=4'b1010;//ʵʱ��ʾʱ��
    #100000
    sw[3:0]=4'b0010;//ʵʱ��ʾʱ��
    #100000
    sw[3:0]=4'b1110;//ʵʱ��ʾ����
    #100000
    sw[3:0]=4'b1010;//ʵʱ��ʾʱ��
    
    #100000
    sw[3:0]=4'b1101;//���������յ�����
    #100000
    key[1:0]=2'b01;//���ǧλ��һ
    #10000000
    key[1:0]=2'b11;
    sw[3:0]=4'b1111;//����ʱ���������
    #100000
    key[1:0]=2'b01;//Сʱ��һ
    #10000000
    key[1:0]=2'b11;  
    #100000
    key[1:0]=2'b01;//Сʱ��һ
    #10000000
    key[1:0]=2'b11;
    #100000
    key[1:0]=2'b10;//���ӵ�����
    #10000000
    key[1:0]=2'b11;  
    #100000
    key[1:0]=2'b01;//���Ӽ�һ
    #10000000
    key[1:0]=2'b11; 
 
    #100000  
    sw[3:0]=4'b1010;//ʵʱ��ʾʱ��
    #10000000
    sw[3:0]=4'b0010;//�ر�����


//    #100000
//    key[1:0]=2'b10;//״̬��ת
//    #100000
    
//        #100000
//    key[1:0]=2'b01;


end
always      begin
#5
    clk_in_p=~clk_in_p;
    clk_in_n=~clk_in_n;
end
endmodule
